library verilog;
use verilog.vl_types.all;
entity SubBytes_TB is
end SubBytes_TB;
