library verilog;
use verilog.vl_types.all;
entity SubBytesLP_TB is
end SubBytesLP_TB;
